module Instruction_Mem(
	input wire [6:0] addr,
	output wire [31:0] data );

//parameter NMEM = 128;   // Number of memory entries, not the same as the memory size
//parameter IM_DATA = "im_data.txt";  // file to read data from
reg [31:0] mem [0:127];  // 32-bit memory with 128 entries

initial
begin
/*
	mem[0] = 32'b100011_00000_10000_00000_00000_000000; // lw s0 0($zero) , s0 = 0 
	mem[1] = 32'b100011_00000_10001_00000_00000_000100; // lw s1 4($zero) , s1 = 0
	mem[2] = 32'b000000_10000_10001_10000_00000_100000; // add s0 s0 s1 , s0 = 0 
	*/

	// $readmemh(IM_DATA, mem, 0, NMEM-1);
	mem[0] = 32'b100011_00000_10000_00000_00000_000000; // lw s0 0($zero) , s0 = 1 
	mem[1] = 32'b100011_00000_10001_00000_00000_000100; // lw s1 4($zero) , s1 = 0
	mem[2] = 32'b000000_10000_10001_10010_00000_100000; // add s2 s0 s1 , s2 = 1 
	mem[3] = 32'b000000_10000_10001_10011_00000_100010; // sub s3 s0 s1 , s3 = 1
	mem[4] = 32'b000000_10010_10011_10100_00000_100100; // and s4 s2 s3 , s4 = 1
	mem[5] = 32'b000000_10010_10011_10101_00000_100110; // xor s5 s2 s3 , s5 = 0
	mem[6] = 32'b000000_10101_10100_10110_00000_101010; // slt s6 s5 s4 , s6 = 1
 	mem[7] = 32'b000100_10101_10001_00000_00000_000001; // beq s5 s1 1 , s5 = s1 = 0
	mem[8] = 32'b000010_00000_00000_00000_00000_001101; // j 13 , it is not executed at first, but is executed after the jump. (mem[12])
	mem[9] = 32'b100011_00000_10111_00000_00000_001000; // lw s7 8($zero) , s7 = 0
	mem[10]= 32'b101011_10111_10101_00000_00000_010000; // sw s5 16(s7) , mem[4] = 0
	mem[11]= 32'b100011_10111_10000_00000_00000_010000; // lw s0 16(s7) , s0 = mem[4] = 0
	mem[12]= 32'b000010_00000_00000_00000_00000_000011; // j 3
	mem[13]= 32'b000000_10000_00000_10111_00000_100111; // nor s7 s0 $zero , s7 = 32'b1111_1111_1111_1111_1111_1111_1111_1111;
	mem[14]= 32'b100011_00000_01000_00000_00000_101000; // lw t0 40($zero) , t0 = 32'b0101_0101_1010_1010_0101_0101_1010_1010;
	mem[15]= 32'b100011_00000_01001_00000_00000_101100; // lw t1 44($zero) , t1 = 32'b0111_0111_1000_1000_0111_0111_1000_1000;
	mem[16]= 32'b000000_01000_01001_01010_00000_100000; // add t2 t0 t1    , t2 = 32'b1100_1101_0011_0010_1100_1101_0011_0010; positive value (overflow)
	mem[17]= 32'b000000_01000_01001_01011_00000_100010; // sub t3 t0 t1    , t3 = 32'b1101_1110_0010_0001_1101_1110_0010_0010; negative value
	mem[18]= 32'b000000_01000_01001_01100_00000_100100; // and t4 t0 t1    , t4 = 32'b0101_0101_1000_1000_0101_0101_1000_1000;
	mem[19]= 32'b000000_01000_01001_01101_00000_100110; // xor t5 t0 t1    , t5 = 32'b0010_0010_0010_0010_0010_0010_0010_0010;
	mem[20]= 32'b000000_01010_01011_01110_00000_101010; // slt t6 t2 t3    , t6 = 32'd1;
	
end

assign data = mem[addr][31:0];

endmodule
